/* VGA Adapter
 *
 * This is a simulated VGA adapter for DESim, which (optionally) includes a video memory. 
 * If the video memory is included, then the VGA controller first draws the contents of this 
 * memory as a background image. Then, it sets the VGA_SYNC signal to indicate that the 
 * VGA controller is in drawing mode. In this mode the controller draws individual pixels 
 * as selected by color, (x,y), write.
 *
 * Three resolutions are supported: 640x480, 320x240, and 160x120. The resolution used should 
 * match whatever is set in the DESim GUI.
*/

module vga_adapter(
            resetn,
            clock,
            color,
            x, y, write,
            VGA_X, 
            VGA_Y, 
            VGA_COLOR, 
            VGA_SYNC,
            plot);
 
    input wire resetn;
    input wire clock;

    // The VGA resolution, which can be set to "640x480", "320x240", and "160x120"
    parameter RESOLUTION = "160x120";
    /* The number of bits used to represent a pixel. An equal number of bits is allocated for 
     * the red (R), green (G) and blue (B) components. Thus, for COLOR_DEPTH = 3, there is one bit
     * for each of the R, G, B components, and eight different colors can be displayed. */
    parameter COLOR_DEPTH = 3;  // default

    input wire [COLOR_DEPTH-1:0] color;

    // Number of VGA pixel X coordinate (column) and Y coordinate (row) bits
    parameter nX = (RESOLUTION == "640x480") ? 10 : ((RESOLUTION == "320x240") ? 9 : 8);
    parameter nY = (RESOLUTION == "640x480") ? 9 : ((RESOLUTION == "320x240") ? 8 : 7);

    parameter BACKGROUND_IMAGE = "background.mif";
    
    input wire [nX-1:0] x;        // used to write to pixels in drawing mode
    input wire [nY-1:0] y;        // used to write to pixels in drawing mode
    input wire write;             // used to write to pixels in drawing mode
    output wire [nX-1:0] VGA_X;   // DESim VGA output
    output wire [nY-1:0] VGA_Y;   // DESim VGA output
    output wire [23:0] VGA_COLOR; // DESim VGA output
    output wire VGA_SYNC;         // set to 1 when in drawing mode
    output wire plot;             // DESim VGA plot output

`ifdef VGA_MEMORY
    // Number of address bits on the video memory
    parameter Mn = (RESOLUTION == "640x480") ? 19 : ((RESOLUTION == "320x240") ? 17 : 15);

    // Number of columns and rows in the video memory
    parameter COLS = (RESOLUTION == "640x480") ? 640 : ((RESOLUTION == "320x240") ? 320 : 160);
    parameter ROWS = (RESOLUTION == "640x480") ? 480 : ((RESOLUTION == "320x240") ? 240 : 120);

    wire [Mn-1:0] controller_to_video_memory_addr; // memory addresses generated by controller
    wire [COLOR_DEPTH-1:0] to_ctrl_color;          // pixel color read from memory

    wire [nX-1:0] VGA_x;                           // needed to support drawing mode
    wire [nY-1:0] VGA_y;                           // needed to support drawing mode
    wire [23:0] VGA_color, color_24;               // needed to support drawing mode
    wire ctrl_plot, VGA_plot, VGA_sync;            // needed to support drawing mode

    /* Create the video memory. This memory is used only to display the background MIF image.
     * This memory is not updated, or used at all, after the MIF has been displayed */
	altsyncram	VideoMemory (
				.address_a (controller_to_video_memory_addr),
				.clock0 (clock),
				.q_a (to_ctrl_color),
				.aclr0 (1'b0),
				.aclr1 (1'b0),
				.address_b (1'b1),
				.addressstall_a (1'b0),
				.addressstall_b (1'b0),
				.byteena_a (1'b1),
				.byteena_b (1'b1),
				.clock1 (1'b1),
				.clocken0 (1'b1),
				.clocken1 (1'b1),
				.clocken2 (1'b1),
				.clocken3 (1'b1),
				.data_a ({COLOR_DEPTH{1'b1}}),
				.data_b (1'b1),
				.eccstatus (),
				.q_b (),
				.rden_a (1'b1),
				.rden_b (1'b1),
				.wren_a (1'b0),
				.wren_b (1'b0));
	defparam
		VideoMemory.address_aclr_a = "NONE",
		VideoMemory.clock_enable_input_a = "BYPASS",
		VideoMemory.clock_enable_output_a = "BYPASS",
		VideoMemory.init_file = "BACKGROUND_IMAGE.mif",
		VideoMemory.intended_device_family = "Cyclone V",
		VideoMemory.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
		VideoMemory.lpm_type = "altsyncram",
		VideoMemory.numwords_a = COLS * ROWS,
		VideoMemory.operation_mode = "ROM",
		VideoMemory.outdata_aclr_a = "NONE",
		VideoMemory.outdata_reg_a = "UNREGISTERED",
		VideoMemory.widthad_a = Mn,
		VideoMemory.width_a = COLOR_DEPTH,
		VideoMemory.width_byteena_a = 1,
        VideoMemory.power_up_uninitialized = "FALSE",
        VideoMemory.init_file = BACKGROUND_IMAGE;

    vga_controller controller(
        .vga_clock(clock),
        .resetn(resetn),
        .pixel_color(to_ctrl_color), // a pixel color from the MIF background
        .memory_address(controller_to_video_memory_addr), // used to read MIF background
        .VGA_X(VGA_x),          // for DESim VGA display
        .VGA_Y(VGA_y),          // for DESim VGA display
        .VGA_COLOR(VGA_color),  // for DESim VGA display
        .VGA_SYNC(VGA_sync),
        .plot(VGA_plot));
        defparam controller.COLOR_DEPTH  = COLOR_DEPTH ;
        defparam controller.nX = nX;
        defparam controller.nY = nY;
        defparam controller.Mn = Mn;
        defparam controller.ROWS = ROWS;
        defparam controller.COLS = COLS;

    // delay sync by one cycle to draw the last pixel of MIF background
    vga_ff USYNC (VGA_sync, resetn, clock, VGA_SYNC);
    /* Before VGA_SYNC becomes 1, draw the background (via the controller).
       But after VGA_SYNC becomes 1, draw pixels using x, y, color, write */
    assign VGA_X = !VGA_SYNC ? VGA_x : x;
    assign VGA_Y = !VGA_SYNC ? VGA_y : y;
    // for color, which is COLOR_DEPTH bits, convert to 24-bit color
    vga_convert UC (color, color_24);
        defparam UC.COLOR_DEPTH = COLOR_DEPTH;
    assign VGA_COLOR = !VGA_SYNC ? VGA_color : color_24; 
    assign plot = !VGA_SYNC ? VGA_plot : write;

`else   // no video memory 

    assign VGA_X = x;
    assign VGA_Y = y;
    vga_convert UC (color, VGA_COLOR);
        defparam UC.COLOR_DEPTH = COLOR_DEPTH;
    assign VGA_SYNC = 1'b1;
    assign plot = write;

`endif // USE_MEMORY

endmodule

// D flip-flop with reset
module vga_ff(D, Resetn, Clock, Q);
    input wire D;
    input wire Resetn, Clock;
    output reg Q;

    always @(posedge Clock)
        if (!Resetn)
            Q <= 1'b0;
        else
            Q <= D;
endmodule

/* Convert COLOR_DEPTH to 24-bit color. The RGB components of color_in are replicated through 
 * the 8-bit RGB components of color_out. For example, if BITS_PER_RGB is 2 and the R 
 * component is R = 2'b10, then the VGA_R component of color_out will be set to 8'b10101010.
*/
module vga_convert(color_in, color_out);
    parameter COLOR_DEPTH = 3;
    parameter BITS_PER_RGB = COLOR_DEPTH / 3;  // default

    input wire [COLOR_DEPTH-1:0] color_in;
    output wire [23:0] color_out;

	integer index;
	integer sub_index;
    reg [7:0] VGA_R, VGA_G, VGA_B;
    always @(*)
	begin		
		VGA_R <= 'b0;
		VGA_G <= 'b0;
		VGA_B <= 'b0;
		for (index = 8-BITS_PER_RGB; index >= 0; index = index - BITS_PER_RGB)
		begin
            for (sub_index = BITS_PER_RGB - 1; sub_index >= 0; sub_index = sub_index - 1)
            begin
                VGA_R[sub_index+index] <= color_in[sub_index + BITS_PER_RGB*2];
                VGA_G[sub_index+index] <= color_in[sub_index + BITS_PER_RGB];
                VGA_B[sub_index+index] <= color_in[sub_index];
            end
        end	
    end
    assign color_out = {VGA_R,VGA_G,VGA_B};

endmodule
